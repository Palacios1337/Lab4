module Status();

endmodule
